-- Dump

/*
 * Copyright 2017, Data61, CSIRO (ABN 41 687 119 230)
 *
 * SPDX-License-Identifier: BSD-2-Clause
 */

arch arm11

objects {

untyped@0xf0000000@12 = ut (12 bits)
untyped@0xf0001000@12 = ut (12 bits)
untyped@0xf0002000@12 = ut (12 bits)
untyped@0xf0003000@12 = ut (12 bits)
untyped@0xf0004000@12 = ut (12 bits)
untyped@0xf0005000@12 = ut (12 bits)
untyped@0xf0006000@12 = ut (12 bits)
untyped@0xf0007000@12 = ut (12 bits)
untyped@0xf0008000@12 = ut (12 bits)
untyped@0xf0009000@12 = ut (12 bits)
untyped@0xf000a000@12 = ut (12 bits)
untyped@0xf000b000@12 = ut (12 bits)
untyped@0xf000c000@12 = ut (12 bits)
untyped@0xf000d000@12 = ut (12 bits)
untyped@0xf000e000@12 = ut (12 bits)
untyped@0xf000f000@12 = ut (12 bits)
untyped@0xf0031800@11 = ut (11 bits)
untyped@0xf0032000@13 = ut (13 bits)
untyped@0xf0034000@14 = ut (14 bits)
untyped@0xf0038000@15 = ut (15 bits)
untyped@0xf0040000@18 = ut (18 bits)
untyped@0xf0080000@19 = ut (19 bits)
untyped@0xf0100000@20 = ut (20 bits)
untyped@0xf0200000@20 = ut (20 bits)
untyped@0xf0300000@14 = ut (14 bits)
untyped@0xf0304000@13 = ut (13 bits)
untyped@0xf0317000@12 = ut (12 bits)
untyped@0xf0318000@15 = ut (15 bits)
untyped@0xf0320000@17 = ut (17 bits)
untyped@0xf0340000@18 = ut (18 bits)
untyped@0xf0380000@19 = ut (19 bits)
untyped@0xf0400000@22 = ut (22 bits)
untyped@0xf0800000@23 = ut (23 bits)
untyped@0xf1000000@24 = ut (24 bits)
untyped@0xf2000000@25 = ut (25 bits)
untyped@0xf4000000@25 = ut (25 bits)
untyped@0xf6000000@24 = ut (24 bits)
untyped@0xf7000000@23 = ut (23 bits)
untyped@0xf7800000@22 = ut (22 bits)
untyped@0xf7c00000@21 = ut (21 bits)
untyped@0xf7e00000@20 = ut (20 bits)
untyped@0xf7f00000@19 = ut (19 bits)
untyped@0xf7f80000@18 = ut (18 bits)
untyped@0xf7fc0000@17 = ut (17 bits)
untyped@0xf7fe0000@15 = ut (15 bits)
untyped@0xf7fe8000@14 = ut (14 bits)
cnode@0xf7ff0000 = cnode(12 bits)
tcb@0xf0031700 = tcb
frame@0x10000000 = frame(1M)
frame@0x10100000 = frame(1M)
frame@0x10200000 = frame(1M)
frame@0x10300000 = frame(1M)
frame@0x10400000 = frame(1M)
frame@0x10500000 = frame(1M)
frame@0x10600000 = frame(1M)
frame@0x10700000 = frame(1M)
frame@0x10800000 = frame(1M)
frame@0x10900000 = frame(1M)
frame@0x10a00000 = frame(1M)
frame@0x10b00000 = frame(1M)
frame@0x10c00000 = frame(1M)
frame@0x10d00000 = frame(1M)
frame@0x10e00000 = frame(1M)
frame@0x10f00000 = frame(1M)
frame@0x11000000 = frame(1M)
frame@0x11100000 = frame(1M)
frame@0x11200000 = frame(1M)
frame@0x11300000 = frame(1M)
frame@0x11400000 = frame(1M)
frame@0x11500000 = frame(1M)
frame@0x11600000 = frame(1M)
frame@0x11700000 = frame(1M)
frame@0x11800000 = frame(1M)
frame@0x11900000 = frame(1M)
frame@0x11a00000 = frame(1M)
frame@0x11b00000 = frame(1M)
frame@0x11c00000 = frame(1M)
frame@0x11d00000 = frame(1M)
frame@0x11e00000 = frame(1M)
frame@0x11f00000 = frame(1M)
frame@0x12000000 = frame(1M)
frame@0x12100000 = frame(1M)
frame@0x12200000 = frame(1M)
frame@0x12300000 = frame(1M)
frame@0x12400000 = frame(1M)
frame@0x12500000 = frame(1M)
frame@0x12600000 = frame(1M)
frame@0x12700000 = frame(1M)
frame@0x12800000 = frame(1M)
frame@0x12900000 = frame(1M)
frame@0x12a00000 = frame(1M)
frame@0x12b00000 = frame(1M)
frame@0x12c00000 = frame(1M)
frame@0x12d00000 = frame(1M)
frame@0x12e00000 = frame(1M)
frame@0x12f00000 = frame(1M)
frame@0x13000000 = frame(1M)
frame@0x13100000 = frame(1M)
frame@0x13200000 = frame(1M)
frame@0x13300000 = frame(1M)
frame@0x13400000 = frame(1M)
frame@0x13500000 = frame(1M)
frame@0x13600000 = frame(1M)
frame@0x13700000 = frame(1M)
frame@0x13800000 = frame(1M)
frame@0x13900000 = frame(1M)
frame@0x13a00000 = frame(1M)
frame@0x13b00000 = frame(1M)
frame@0x13c00000 = frame(1M)
frame@0x13d00000 = frame(1M)
frame@0x13e00000 = frame(1M)
frame@0x13f00000 = frame(1M)
frame@0x18000000 = frame(1M)
frame@0x18100000 = frame(1M)
frame@0x18200000 = frame(1M)
frame@0x18300000 = frame(1M)
frame@0x18400000 = frame(1M)
frame@0x18500000 = frame(1M)
frame@0x18600000 = frame(1M)
frame@0x18700000 = frame(1M)
frame@0x18800000 = frame(1M)
frame@0x18900000 = frame(1M)
frame@0x18a00000 = frame(1M)
frame@0x18b00000 = frame(1M)
frame@0x18c00000 = frame(1M)
frame@0x18d00000 = frame(1M)
frame@0x18e00000 = frame(1M)
frame@0x18f00000 = frame(1M)
frame@0x19000000 = frame(1M)
frame@0x19100000 = frame(1M)
frame@0x19200000 = frame(1M)
frame@0x19300000 = frame(1M)
frame@0x19400000 = frame(1M)
frame@0x19500000 = frame(1M)
frame@0x19600000 = frame(1M)
frame@0x19700000 = frame(1M)
frame@0x19800000 = frame(1M)
frame@0x19900000 = frame(1M)
frame@0x19a00000 = frame(1M)
frame@0x19b00000 = frame(1M)
frame@0x19c00000 = frame(1M)
frame@0x19d00000 = frame(1M)
frame@0x19e00000 = frame(1M)
frame@0x19f00000 = frame(1M)
frame@0x30000000 = frame(1M)
frame@0x30100000 = frame(1M)
frame@0x30200000 = frame(1M)
frame@0x30300000 = frame(1M)
frame@0x30400000 = frame(1M)
frame@0x30500000 = frame(1M)
frame@0x30600000 = frame(1M)
frame@0x30700000 = frame(1M)
frame@0x30800000 = frame(1M)
frame@0x30900000 = frame(1M)
frame@0x30a00000 = frame(1M)
frame@0x30b00000 = frame(1M)
frame@0x30c00000 = frame(1M)
frame@0x30d00000 = frame(1M)
frame@0x30e00000 = frame(1M)
frame@0x30f00000 = frame(1M)
frame@0x31000000 = frame(1M)
frame@0x31100000 = frame(1M)
frame@0x31200000 = frame(1M)
frame@0x31300000 = frame(1M)
frame@0x31400000 = frame(1M)
frame@0x31500000 = frame(1M)
frame@0x31600000 = frame(1M)
frame@0x31700000 = frame(1M)
frame@0x31800000 = frame(1M)
frame@0x31900000 = frame(1M)
frame@0x31a00000 = frame(1M)
frame@0x31b00000 = frame(1M)
frame@0x31c00000 = frame(1M)
frame@0x31d00000 = frame(1M)
frame@0x31e00000 = frame(1M)
frame@0x31f00000 = frame(1M)
frame@0x26000000 = frame(4k)
frame@0xb3f80000 = frame(4k)
frame@0xb3f84000 = frame(4k)
frame@0xb3f88000 = frame(4k)
frame@0xb3f8c000 = frame(4k)
frame@0xb3f94000 = frame(4k)
frame@0xb3f98000 = frame(4k)
frame@0xb3f9c000 = frame(4k)
frame@0xb3fa0000 = frame(4k)
frame@0xb3fa4000 = frame(4k)
frame@0xb3fa8000 = frame(4k)
frame@0xb3fac000 = frame(4k)
frame@0xb3fb0000 = frame(4k)
frame@0xb3fb4000 = frame(4k)
frame@0xc0004000 = frame(4k)
frame@0xc0008000 = frame(4k)
frame@0xc000c000 = frame(4k)
frame@0xc0010000 = frame(4k)
frame@0xc0014000 = frame(4k)
frame@0xc0018000 = frame(4k)
frame@0xc001c000 = frame(4k)
frame@0xc0020000 = frame(4k)
frame@0xc0024000 = frame(4k)
frame@0xc0028000 = frame(4k)
frame@0xc003c000 = frame(4k)
frame@0xc3f80000 = frame(4k)
frame@0xc3f84000 = frame(4k)
frame@0xc3f8c000 = frame(4k)
frame@0xc3f90000 = frame(4k)
frame@0xc3f98000 = frame(4k)
frame@0xc3fa4000 = frame(4k)
frame@0xc3fb0000 = frame(4k)
frame@0xc3fc4000 = frame(4k)
frame@0xc3fcc000 = frame(4k)
frame@0xc3fd0000 = frame(4k)
frame@0xc3fd8000 = frame(4k)
frame@0xc3fe0000 = frame(4k)
frame@0xc3fec000 = frame(4k)
frame@0xf002f000 = frame(4k)
frame@0xf0030000 = frame(4k)
frame@0xf0307000 = frame(4k)
frame@0xf0308000 = frame(4k)
frame@0xf0309000 = frame(4k)
frame@0xf030a000 = frame(4k)
frame@0xf030b000 = frame(4k)
frame@0xf030c000 = frame(4k)
frame@0xf030d000 = frame(4k)
frame@0xf030e000 = frame(4k)
frame@0xf030f000 = frame(4k)
frame@0xf0310000 = frame(4k)
frame@0xf0311000 = frame(4k)
frame@0xf0312000 = frame(4k)
frame@0xf0313000 = frame(4k)
frame@0xf0314000 = frame(4k)
frame@0xf0315000 = frame(4k)
frame@0xf0316000 = frame(4k)
pt@0xf0031000 = pt
pd@0xf7fec000 = pd
asid_pool@0xf0306000 = asid_pool (asid_high: 0x0)

} caps {

tcb@0xf0031700{
  0x0: cnode@0xf7ff0000 (guard:0x0, guard_size: 20)
  0x1: pd@0xf7fec000 (asid: (0x0, 0x1))
  0x2: tcb@0xf0031700 (master_reply)
  0x4: frame@0xf002f000 (RW, asid: (0x0, 0x1))
}
cnode@0xf7ff0000{
  0x1: tcb@0xf0031700
  0x2: cnode@0xf7ff0000 (guard:0x0, guard_size: 20)
  0x3: pd@0xf7fec000 (asid: (0x0, 0x1))
  0x4: irq_control
  0x5: asid_control
  0x6: asid_pool@0xf0306000
  0x9: frame@0xf0030000 (RW, asid: (0x0, 0x1))
  0xa: frame@0xf002f000 (RW, asid: (0x0, 0x1))
  0xb: frame@0xf0307000 (RW, asid: (0x0, 0x1))
  0xc: frame@0xf0308000 (RW, asid: (0x0, 0x1))
  0xd: frame@0xf0309000 (RW, asid: (0x0, 0x1))
  0xe: frame@0xf030a000 (RW, asid: (0x0, 0x1))
  0xf: frame@0xf030b000 (RW, asid: (0x0, 0x1))
  0x10: frame@0xf030c000 (RW, asid: (0x0, 0x1))
  0x11: frame@0xf030d000 (RW, asid: (0x0, 0x1))
  0x12: frame@0xf030e000 (RW, asid: (0x0, 0x1))
  0x13: frame@0xf030f000 (RW, asid: (0x0, 0x1))
  0x14: frame@0xf0310000 (RW, asid: (0x0, 0x1))
  0x15: frame@0xf0311000 (RW, asid: (0x0, 0x1))
  0x16: frame@0xf0312000 (RW, asid: (0x0, 0x1))
  0x17: frame@0xf0313000 (RW, asid: (0x0, 0x1))
  0x18: frame@0xf0314000 (RW, asid: (0x0, 0x1))
  0x19: frame@0xf0315000 (RW, asid: (0x0, 0x1))
  0x1a: frame@0xf0316000 (RW, asid: (0x0, 0x1))
  0x1b: pt@0xf0031000 (asid: (0x0, 0x1))
  0x1c: untyped@0xf0000000@12
  0x1d: untyped@0xf0001000@12
  0x1e: untyped@0xf0002000@12
  0x1f: untyped@0xf0003000@12
  0x20: untyped@0xf0004000@12
  0x21: untyped@0xf0005000@12
  0x22: untyped@0xf0006000@12
  0x23: untyped@0xf0007000@12
  0x24: untyped@0xf0008000@12
  0x25: untyped@0xf0009000@12
  0x26: untyped@0xf000a000@12
  0x27: untyped@0xf000b000@12
  0x28: untyped@0xf000c000@12
  0x29: untyped@0xf000d000@12
  0x2a: untyped@0xf000e000@12
  0x2b: untyped@0xf000f000@12
  0x2c: untyped@0xf0031800@11
  0x2d: untyped@0xf0032000@13
  0x2e: untyped@0xf0304000@13
  0x2f: untyped@0xf0034000@14
  0x30: untyped@0xf0300000@14
  0x31: untyped@0xf0038000@15
  0x32: untyped@0xf0040000@18
  0x33: untyped@0xf0080000@19
  0x34: untyped@0xf0100000@20
  0x35: untyped@0xf0200000@20
  0x36: untyped@0xf0317000@12
  0x37: untyped@0xf7fe8000@14
  0x38: untyped@0xf0318000@15
  0x39: untyped@0xf7fe0000@15
  0x3a: untyped@0xf0320000@17
  0x3b: untyped@0xf7fc0000@17
  0x3c: untyped@0xf0340000@18
  0x3d: untyped@0xf7f80000@18
  0x3e: untyped@0xf0380000@19
  0x3f: untyped@0xf7f00000@19
  0x40: untyped@0xf7e00000@20
  0x41: untyped@0xf7c00000@21
  0x42: untyped@0xf0400000@22
  0x43: untyped@0xf7800000@22
  0x44: untyped@0xf0800000@23
  0x45: untyped@0xf7000000@23
  0x46: untyped@0xf1000000@24
  0x47: untyped@0xf6000000@24
  0x48: untyped@0xf2000000@25
  0x49: untyped@0xf4000000@25
  0x4a: frame@0xb3f80000 (RW)
  0x4b: frame@0xb3f84000 (RW)
  0x4c: frame@0xb3f88000 (RW)
  0x4d: frame@0xb3f8c000 (RW)
  0x4e: frame@0xb3f94000 (RW)
  0x4f: frame@0xb3f98000 (RW)
  0x50: frame@0xb3f9c000 (RW)
  0x51: frame@0xb3fa0000 (RW)
  0x52: frame@0xb3fa4000 (RW)
  0x53: frame@0xb3fa8000 (RW)
  0x54: frame@0xb3fac000 (RW)
  0x55: frame@0xb3fb0000 (RW)
  0x56: frame@0xb3fb4000 (RW)
  0x57: frame@0xc0004000 (RW)
  0x58: frame@0xc0008000 (RW)
  0x59: frame@0xc000c000 (RW)
  0x5a: frame@0xc0010000 (RW)
  0x5b: frame@0xc0014000 (RW)
  0x5c: frame@0xc0018000 (RW)
  0x5d: frame@0xc001c000 (RW)
  0x5e: frame@0xc0020000 (RW)
  0x5f: frame@0xc0024000 (RW)
  0x60: frame@0xc0028000 (RW)
  0x61: frame@0xc003c000 (RW)
  0x62: frame@0xc3f80000 (RW)
  0x63: frame@0xc3f84000 (RW)
  0x64: frame@0xc3f8c000 (RW)
  0x65: frame@0xc3f90000 (RW)
  0x66: frame@0xc3f98000 (RW)
  0x67: frame@0xc3fa4000 (RW)
  0x68: frame@0xc3fb0000 (RW)
  0x69: frame@0xc3fc4000 (RW)
  0x6a: frame@0xc3fcc000 (RW)
  0x6b: frame@0xc3fd0000 (RW)
  0x6c: frame@0xc3fd8000 (RW)
  0x6d: frame@0xc3fe0000 (RW)
  0x6e: frame@0xc3fec000 (RW)
  0x6f: frame@0x10000000 (RW)
  0x70: frame@0x10100000 (RW)
  0x71: frame@0x10200000 (RW)
  0x72: frame@0x10300000 (RW)
  0x73: frame@0x10400000 (RW)
  0x74: frame@0x10500000 (RW)
  0x75: frame@0x10600000 (RW)
  0x76: frame@0x10700000 (RW)
  0x77: frame@0x10800000 (RW)
  0x78: frame@0x10900000 (RW)
  0x79: frame@0x10a00000 (RW)
  0x7a: frame@0x10b00000 (RW)
  0x7b: frame@0x10c00000 (RW)
  0x7c: frame@0x10d00000 (RW)
  0x7d: frame@0x10e00000 (RW)
  0x7e: frame@0x10f00000 (RW)
  0x7f: frame@0x11000000 (RW)
  0x80: frame@0x11100000 (RW)
  0x81: frame@0x11200000 (RW)
  0x82: frame@0x11300000 (RW)
  0x83: frame@0x11400000 (RW)
  0x84: frame@0x11500000 (RW)
  0x85: frame@0x11600000 (RW)
  0x86: frame@0x11700000 (RW)
  0x87: frame@0x11800000 (RW)
  0x88: frame@0x11900000 (RW)
  0x89: frame@0x11a00000 (RW)
  0x8a: frame@0x11b00000 (RW)
  0x8b: frame@0x11c00000 (RW)
  0x8c: frame@0x11d00000 (RW)
  0x8d: frame@0x11e00000 (RW)
  0x8e: frame@0x11f00000 (RW)
  0x8f: frame@0x12000000 (RW)
  0x90: frame@0x12100000 (RW)
  0x91: frame@0x12200000 (RW)
  0x92: frame@0x12300000 (RW)
  0x93: frame@0x12400000 (RW)
  0x94: frame@0x12500000 (RW)
  0x95: frame@0x12600000 (RW)
  0x96: frame@0x12700000 (RW)
  0x97: frame@0x12800000 (RW)
  0x98: frame@0x12900000 (RW)
  0x99: frame@0x12a00000 (RW)
  0x9a: frame@0x12b00000 (RW)
  0x9b: frame@0x12c00000 (RW)
  0x9c: frame@0x12d00000 (RW)
  0x9d: frame@0x12e00000 (RW)
  0x9e: frame@0x12f00000 (RW)
  0x9f: frame@0x13000000 (RW)
  0xa0: frame@0x13100000 (RW)
  0xa1: frame@0x13200000 (RW)
  0xa2: frame@0x13300000 (RW)
  0xa3: frame@0x13400000 (RW)
  0xa4: frame@0x13500000 (RW)
  0xa5: frame@0x13600000 (RW)
  0xa6: frame@0x13700000 (RW)
  0xa7: frame@0x13800000 (RW)
  0xa8: frame@0x13900000 (RW)
  0xa9: frame@0x13a00000 (RW)
  0xaa: frame@0x13b00000 (RW)
  0xab: frame@0x13c00000 (RW)
  0xac: frame@0x13d00000 (RW)
  0xad: frame@0x13e00000 (RW)
  0xae: frame@0x13f00000 (RW)
  0xaf: frame@0x18000000 (RW)
  0xb0: frame@0x18100000 (RW)
  0xb1: frame@0x18200000 (RW)
  0xb2: frame@0x18300000 (RW)
  0xb3: frame@0x18400000 (RW)
  0xb4: frame@0x18500000 (RW)
  0xb5: frame@0x18600000 (RW)
  0xb6: frame@0x18700000 (RW)
  0xb7: frame@0x18800000 (RW)
  0xb8: frame@0x18900000 (RW)
  0xb9: frame@0x18a00000 (RW)
  0xba: frame@0x18b00000 (RW)
  0xbb: frame@0x18c00000 (RW)
  0xbc: frame@0x18d00000 (RW)
  0xbd: frame@0x18e00000 (RW)
  0xbe: frame@0x18f00000 (RW)
  0xbf: frame@0x19000000 (RW)
  0xc0: frame@0x19100000 (RW)
  0xc1: frame@0x19200000 (RW)
  0xc2: frame@0x19300000 (RW)
  0xc3: frame@0x19400000 (RW)
  0xc4: frame@0x19500000 (RW)
  0xc5: frame@0x19600000 (RW)
  0xc6: frame@0x19700000 (RW)
  0xc7: frame@0x19800000 (RW)
  0xc8: frame@0x19900000 (RW)
  0xc9: frame@0x19a00000 (RW)
  0xca: frame@0x19b00000 (RW)
  0xcb: frame@0x19c00000 (RW)
  0xcc: frame@0x19d00000 (RW)
  0xcd: frame@0x19e00000 (RW)
  0xce: frame@0x19f00000 (RW)
  0xcf: frame@0x26000000 (RW)
  0xd0: frame@0x30000000 (RW)
  0xd1: frame@0x30100000 (RW)
  0xd2: frame@0x30200000 (RW)
  0xd3: frame@0x30300000 (RW)
  0xd4: frame@0x30400000 (RW)
  0xd5: frame@0x30500000 (RW)
  0xd6: frame@0x30600000 (RW)
  0xd7: frame@0x30700000 (RW)
  0xd8: frame@0x30800000 (RW)
  0xd9: frame@0x30900000 (RW)
  0xda: frame@0x30a00000 (RW)
  0xdb: frame@0x30b00000 (RW)
  0xdc: frame@0x30c00000 (RW)
  0xdd: frame@0x30d00000 (RW)
  0xde: frame@0x30e00000 (RW)
  0xdf: frame@0x30f00000 (RW)
  0xe0: frame@0x31000000 (RW)
  0xe1: frame@0x31100000 (RW)
  0xe2: frame@0x31200000 (RW)
  0xe3: frame@0x31300000 (RW)
  0xe4: frame@0x31400000 (RW)
  0xe5: frame@0x31500000 (RW)
  0xe6: frame@0x31600000 (RW)
  0xe7: frame@0x31700000 (RW)
  0xe8: frame@0x31800000 (RW)
  0xe9: frame@0x31900000 (RW)
  0xea: frame@0x31a00000 (RW)
  0xeb: frame@0x31b00000 (RW)
  0xec: frame@0x31c00000 (RW)
  0xed: frame@0x31d00000 (RW)
  0xee: frame@0x31e00000 (RW)
  0xef: frame@0x31f00000 (RW)
}
pd@0xf7fec000{
  0x0: pt@0xf0031000
}
pt@0xf0031000{
  0x7: frame@0xf0307000 (RW)
  0x8: frame@0xf0308000 (RW)
  0x9: frame@0xf0309000 (RW)
  0xa: frame@0xf030a000 (RW)
  0xb: frame@0xf030b000 (RW)
  0xc: frame@0xf030c000 (RW)
  0xd: frame@0xf030d000 (RW)
  0xe: frame@0xf030e000 (RW)
  0xf: frame@0xf030f000 (RW)
  0x10: frame@0xf0310000 (RW)
  0x11: frame@0xf0311000 (RW)
  0x12: frame@0xf0312000 (RW)
  0x13: frame@0xf0313000 (RW)
  0x14: frame@0xf0314000 (RW)
  0x15: frame@0xf0315000 (RW)
  0x16: frame@0xf0316000 (RW)
  0x17: frame@0xf002f000 (RW)
  0x18: frame@0xf0030000 (RW)
}
asid_pool@0xf0306000{
  0x1: pd@0xf7fec000
}

} cdt {

(cnode@0xf7ff0000,0x2) {(tcb@0xf0031700,0x0)}
(cnode@0xf7ff0000,0x3) {(tcb@0xf0031700,0x1)}
(cnode@0xf7ff0000,0xa) {(tcb@0xf0031700,0x4)}

}
